`define TIMER_CTRL_ADDR  8'h0
`define TIMER_CTRL_IN_ADDR  8'h1
`define TIMER_CTRL_OUT_ADDR  8'h2
`define TIMER_STATUS_ADDR 8'h4
`define TIMER_CNT_INIT_ADDR 8'h8
`define TIMER_CNT_MIN_ADDR 8'h9
`define TIMER_CNT_MAX_ADDR 8'hA
`define TIMER_CNT_ADDR 8'hB
`define TIMER_CNT_MATCH_0_ADDR 8'hC
`define TIMER_CNT_MATCH_1_ADDR 8'hD
