`SHOWM(Input pulses counter);

reg_read(`TIMER_CTRL_ADDR);
//reg_write(`TIMER_CTRL_ADDR,8'h01);
reg_write(`TIMER_CNT_MAX_ADDR,8'd10);
reg_write(`TIMER_CTRL_ADDR,8'h09);
delay(1000);
