
// Блок генерации ШИМ
module PWM_block #(
	parameter	COUNTER_SIZE  = 32,
					NUM_COMP  = 2)
	(
		input logic rst,												// Сброс
		input logic clk,												// Тактирование
		input logic en,												// Разрешение работы
		input logic [NUM_COMP-1:0] [COUNTER_SIZE-1:0] match_value,
		input logic [COUNTER_SIZE-1:0] counter_value,
		input logic [NUM_COMP-1:0] intr_en,
		input logic [NUM_COMP-1:0] trg_en,     
		input logic pwm_mode,										// Режим ШИМ
		input	logic inv,												// Инверсия

		output logic timer_out,trigger,
		output [NUM_COMP-1:0] intr,      
		output logic [NUM_COMP-1:0] match						// Совпадение
		);

reg timer_out_internal;

	wire high_pwm;														// Активный уровень
	wire low_pwm;
	reg [NUM_COMP-1:0] 	match_past;
	wire [NUM_COMP-1:0]	match_rise;
	wire [NUM_COMP-1:0]	trigger_internal;
	logic [NUM_COMP-1:0]	local_match_flag;												// Для организации локальной связи без внешнего модуля
	assign trigger = |trigger_internal;

	// Задаем количество ШИМ каналов.
	// ШИМ работает в классическом режиме. В перспективе можно добавить режим "ШИМ с точной фазой"
	genvar a;
	generate
		for (a = 0; a < NUM_COMP; a=a+1)	begin: interrupt_unit
			assign match[a] = (match_value[a] == counter_value);
			assign match_rise[a] = (~match_past[a] & match[a]);
		end
	 
	for (a = 0;a < NUM_COMP; a=a+1 )	begin: compare_unit
		assign trigger_internal[a] = (match[a] & trg_en[a]);
		end 
		
	endgenerate
	
	always @ (posedge clk or posedge rst) begin
		if (rst)	match_past = 0;
			else	match_past = match;  
	end  


// Блок генерации ШИМ
// устанавливается при совпадении с 0
// не установлен, если комп совпадает с 1

assign high_pwm = match_rise[0] & en & pwm_mode;  
assign low_pwm  = match_rise[1] & en & pwm_mode;

	always @ (posedge clk or posedge rst) begin
	if (rst)	timer_out_internal	=	0;											// При сброре обнуляем интервал
		else	if (high_pwm)	timer_out_internal	=	1;						// 
				else if (low_pwm)	timer_out_internal =	0;
						else 	timer_out_internal = timer_out_internal;    
	end


	
assign local_match_flag = match;
assign intr = (intr_en & local_match_flag );
assign timer_out = inv	?	(~timer_out_internal)	:	(timer_out_internal);

endmodule
