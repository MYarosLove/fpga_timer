`define TB_SCOPE  tb_counter
`define TOP_SCOPE `TB_SCOPE.timer
